module RegisterFile (
    input clk, reset,
    input [4:0] rs_address, rt_address, rd_address,
    input [31:0] rs_data, rt_data,
    input write_enable,
    output reg [31:0] rs_out, rt_out
);



endmodule